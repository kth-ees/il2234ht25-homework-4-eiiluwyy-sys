
module adder16(
  input  logic [15:0] a,
  input  logic [15:0] b,
  output logic [15:0] sum
);
  assign sum = a + b;
endmodule
