
module subtractor16(
  input  logic [15:0] a,
  input  logic [15:0] b,
  output logic [15:0] diff
);
  assign diff = a - b;
endmodule
